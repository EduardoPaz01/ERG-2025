* Symmetric-Source
*
* SPICE MODEL (by EduardoPaz01)
* SUBCIRCUIT
*
* Connections:
.SUBCKT symmetric_source IN+ IN- GND +8V -8V
L1 IN+ IN- 1.713H
L2 N001 0 2.87mH
L3 0 N004 2.87mH
D1 N001 N002 1N4007
D3 N003 N001 1N4007
D4 N004 N002 1N4007
D5 N003 N004 1N4007
X§U1 N002 0 +8V LM7808 ;§pnba IN)GND)OUT
X§U2 N003 0 -8V LM7908 ;§pnba IN)GND)OUT
C4 0 -8V 100nF V=35V
C6 0 -8V 100µ V=25 Irms=145m Rser=0.62 Lser=0 mfg="Nichicon" pn="UPR1E101MPH" type="Al electrolytic"
C2 0 N003 2200µ V=25 Irms=2.39 Rser=0.021 Lser=0 mfg="Panasonic" pn="ECA1EFQ222L" type="Al electrolytic"
C1 N002 0 2200µ V=25 Irms=2.39 Rser=0.021 Lser=0 mfg="Panasonic" pn="ECA1EFQ222L" type="Al electrolytic"
C3 +8V 0 100µ V=25 Irms=145m Rser=0.62 Lser=0 mfg="Nichicon" pn="UPR1E101MPH" type="Al electrolytic"
C5 +8V 0 100nF V=35V
.model D D
.lib C:\Users\Acer\AppData\Local\LTspice\lib\cmp\standard.dio
K L1 L2 L3 1.
.lib C:\Users\Acer\repos\ERG-2025\symmetric-source\SPICE-models\LM7808.CIR
.lib C:\Users\Acer\repos\ERG-2025\symmetric-source\SPICE-models\LM7908.CIR
.ENDS symmetric_source
