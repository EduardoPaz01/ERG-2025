* LM7808
*
* SPICE MODEL (adapted by EduardoPaz01)
* SUBCIRCUIT
*
* Connections: In Gnd Out
.SUBCKT LM7808 IN GND OUT
RBIAS 40 OUT 220
RADJ GND 40 1188
D4 4 OUT D_Z6V0
D3 5 6 D_Z6V3
D2 7 IN D_Z6V3
D1 OUT 8 D_Z6V3
QT26 IN 10 9 Q_NPN 20.0
QT25 IN 11 10 Q_NPN 2.0
QT24_2 13 12 5 Q_NPN 0.1
QT24 13 12 14 Q_NPN 0.1
QT23 17 16 15 Q_NPN 1.0
QT21 19 18 OUT Q_NPN 0.1
QT19 21 OUT 20 Q_NPN 1.0
QT17 23 OUT 22 Q_NPN 0.1
QT13 IN 25 24 Q_NPN 0.1
QT11 16 27 26 Q_NPN 0.1
QT7 30 29 28 Q_NPN 0.1
QT5 29 31 OUT Q_NPN 0.1
QT3 33 31 32 Q_NPN 0.1
QT22_2 17 17 IN Q_PNP 1.0
QT22 16 17 IN Q_PNP 1.0
QT20 OUT 19 16 Q_PNP 0.1
QT18 21 21 16 Q_PNP 0.1
QT16 23 21 16 Q_PNP 0.1
QT15 OUT 23 25 Q_PNP 0.1
QT12 OUT 24 16 Q_PNP 0.1
QT9 27 30 34 Q_PNP 0.1
QT6 OUT 29 34 Q_PNP 0.1
QT14 25 33 35 Q_PNP 0.1
QT10 16 33 36 Q_PNP 0.1
QT8 34 33 37 Q_PNP 0.1
QT4 31 33 38 Q_PNP 0.1
QT2 33 33 39 Q_PNP 0.1
R27 4 40 50
R26 9 OUT 100M
R25 9 14 2
R24 5 14 160
R23 7 6 18K
R22 10 OUT 160
R21 12 13 400
R20 18 13 13K
R19 16 11 370
R18 15 10 130
R17 16 12 12K
C3 19 18 5P
R16 16 19 6.7K
R15 20 22 2.4K
R14 22 4 12K
C2 23 4 30P
C1 23 OUT 30P
R13 24 OUT 5.1K
R12 26 OUT 72
R11 27 OUT 5.8K
R10 28 OUT 4.1K
R9 32 OUT 180
R8 34 30 12.4K
R7 31 29 130
R6 8 31 100K
R5 IN 35 5.6K
R4 IN 36 82
R3 IN 37 190
R2 IN 38 310
R1 IN 39 310
JT1 IN OUT 8 J_N
.MODEL D_Z6V0 D(IS=10F N=1.04 BV=6.0 IBV=1M CJO = 1P TT = 10p)
.MODEL D_Z6V3 D(IS=10F N=1.04 BV=6.3 IBV=1M CJO = 1P TT = 10p)
.MODEL Q_NPN NPN(IS=10F NF=1.04 NR=1.04 BF=100 CJC=1P CJE=2P TF=10P TR=1N VAF=90)
.MODEL Q_PNP PNP(IS=10F NF=1.04 NR=1.04 BF=50 CJC=1P CJE=2P TF=10P TR=1N VAF=45)
.MODEL J_N NJF(VTO=-7)
.ENDS
